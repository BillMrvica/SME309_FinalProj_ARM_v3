`timescale 1ns / 1ps
// The multiplier template is provided, and you should modify it to the improved one and share the hardware resource to implement division.
//�ṩ�˳˷���ģ�壬��Ӧ�ý����޸�Ϊ�Ľ���ģ�壬������Ӳ����Դ��ʵ�ֳ�����
module MCycle
  #(parameter width = 32) // 32-bits for ARMv3
   (
     input CLK,   // Connect to CPU clock
     input Reset, // Connect to the reset of the ARM processor.
     input Start_MCycle, // Multi-cycle Enable. The control unit should assert this when MUL or DIV instruction is detected.
     input MCycleOp_MCycle, // Multi-cycle Operation. "0" for unsigned multiplication, "1" for unsigned division. Generated by Control unit.
     input [width-1:0] Operand1_MCycle, // Multiplicand / Dividend
     input [width-1:0] Operand2_MCycle, // Multiplier / Divisor
     output [width-1:0] Result_MCycle,  //For MUL, assign the lower-32bits result; For DIV, assign the quotient.
     output reg Busy_MCycle // Set immediately when Start_MCycle is set. Cleared when the Results become ready. This bit can be used to stall the processor while multi-cycle operations are on.
   );

  localparam IDLE = 1'b0;
  localparam COMPUTING = 1'b1;
  reg state, n_state;
  reg done;
  // state machine
always @(posedge CLK or posedge Reset)
  begin
    if(Reset)
      state <= IDLE;
    else
      state <= n_state;
  end

always @(*)
  begin
    case(state)
      IDLE:begin
                if(Start_MCycle) begin
                    n_state = COMPUTING;
                    Busy_MCycle = 1'b1;
                end else begin
                    n_state = IDLE;
                    Busy_MCycle = 1'b0;
                end
           end
      COMPUTING:begin
                    if(~done)begin
                        n_state = COMPUTING ;
                        Busy_MCycle = 1'b1 ;
                    end else begin
                        n_state = IDLE;
                        Busy_MCycle = 1'b0;
                    end
                end
    endcase
end

reg [5:0] count = 0 ; // assuming no computation takes more than 64 cycles.����û�м�����Ҫ����64�����ڡ�
reg [2*width:0] temp_sum2 = 0 ;
reg [2*width:0] shifted_op2_divider_mul ;
reg [2*width:0] temp_sum_divider_mul;
  // Multi-cycle Multiplier & divider
always@(posedge CLK or posedge Reset)
  begin: COMPUTING_PROCESS // process which does the actual computation
    if( Reset )
    begin
      count <= 0 ;
      shifted_op2_divider_mul <= {  {1'b0},Operand2_MCycle,{width{1'b0}} } ;
      temp_sum_divider_mul <={  {1'b0},{width{1'b0}} ,Operand1_MCycle};
      done <= 0;
    end
    // state: IDLE
    else if(state == IDLE)
    begin
      if(n_state == COMPUTING)
      begin
        count <= 0 ;
        shifted_op2_divider_mul <= {  {1'b0},Operand2_MCycle,{width{1'b0}} } ;
        temp_sum_divider_mul <={  {1'b0},{width{1'b0}} ,Operand1_MCycle};
        done <= 0;
      end
      // else IDLE->IDLE: registers unchanged
    end
    // state: COMPUTING
    else if(n_state == COMPUTING)
    begin
      if( ~MCycleOp_MCycle )
      begin // Multiply operation
        // The intial version of multiplier template, modify it to the improved one
        if(count == width-1)
        begin // last cycle
          done <= 1'b1 ;
          count <= 0;
        end
        else
        begin
          done <= 1'b0;
          count <= count + 1;
        end
        if(temp_sum_divider_mul[0]) begin
            temp_sum2 = shifted_op2_divider_mul + temp_sum_divider_mul;
            temp_sum_divider_mul <= {1'b0,temp_sum2[2*width-1 : 1] };
          end else begin 
            temp_sum_divider_mul <= {1'b0, temp_sum_divider_mul[2*width-1 : 1]} ;
          end
        // else temp_sum unchanged        
      end
      // Multiplier end
      else
      begin // Divide operation
        //
        // Fit with your code to design divider, remember to share the hardware resource with the improved multiplier
        //
        if(count == width) begin // last cycle
            done <= 1'b1 ;
            count <= 0;
        end else begin
            done <= 1'b0;
            count <= count + 1;
        end
        temp_sum2 = temp_sum_divider_mul - shifted_op2_divider_mul;
        if(temp_sum2[2*width]) begin
            temp_sum_divider_mul <= { temp_sum_divider_mul[2*width-1 : 0],1'b0};
        end else begin
            temp_sum_divider_mul <= { temp_sum2[2*width : 0],1'b1};
        end
      end
    end
  end
    
assign Result_MCycle = temp_sum_divider_mul[width-1:0];

endmodule


